library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

ENTITY kara256bit_tb IS END kara256bit_tb;
architecture test1 of kara256bit_tb is

SIGNAL t_clk: std_logic:='0';
SIGNAL t_start: std_logic;
SIGNAL t_rst:std_logic;
SIGNAL t_multiplier:unsigned(255 downto 0); 
SIGNAL t_multiplicand:unsigned(255 downto 0);
SIGNAL t_p :unsigned(511 downto 0);
SIGNAL t_done: std_logic;
begin
    UUT : entity work.kara256bit PORT MAP(t_clk,t_start,t_rst,t_multiplier,t_multiplicand,t_p,t_done);
    t_clk <= NOT t_clk AFTER 5 ns;
    PROCESS 
    BEGIN
      WAIT FOR 1 ps;
      --t_multiplier <="1000100011111011001101100001101100001110000000101000101101000010110101101010110011111000111010000010001010100000000010010010111100110001110110011010011001011101110101011111010011010000110010000001100000111111101100111001110001001111110111011100010001001111";
      --t_multiplicand <="1101110100110001100100101000000101010011001110010001001101100001010110010101011101100011110011110000010001001011111110111001010000000111010111011001010000101011010000101010010101101010000011111111110010001100001000001100000011001101101001000110000011000110";
      t_multiplier <="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100001111";
      t_multiplicand <="0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101111";
      t_start <='0';
      t_rst <='0';
      WAIT FOR 40 ns;
      t_start <='1';
      WAIT FOR 10 ns;
      t_start <='0';
      WAIT;
  
    END PROCESS;
end test1 ;

-- inp1 = 1000100011111011001101100001101100001110000000101000101101000010110101101010110011111000111010000010001010100000000010010010111100110001110110011010011001011101110101011111010011010000110010000001100000111111101100111001110001001111110111011100010001001111 
-- inp2 = 1101110100110001100100101000000101010011001110010001001101100001010110010101011101100011110011110000010001001011111110111001010000000111010111011001010000101011010000101010010101101010000011111111110010001100001000001100000011001101101001000110000011000110

-- res = 6198858940839361893948978270737012004036340944350875035352817072789619343786243960855029428733021486480529930089876368607594397724657071869830231096259866
-- reshex = 765B642F2E3F8F2D6B6541B1C0A3A562BE808D556C8E89BCF90F7A0AF210A19C65AB3CFC0F3412C003215CCE40AF3A89120F149EE9C57FDB9EC8645DF4BF751A


